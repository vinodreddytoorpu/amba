package amba_environment_package;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import apb5_environment_package::*;

  `include "amba_defines.sv"
  `include "amba_environment_config.sv"
  `include "amba_virtual_sequencer.sv"
  `include "amba_apb5_requester_subscriber.sv"
  `include "amba_environment.sv"

endpackage : amba_environment_package
