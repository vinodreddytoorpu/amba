
`define AMBA_APB5_ADDR_WIDTH      32
`define AMBA_APB5_DATA_WIDTH      32
`define AMBA_APB5_USER_REQ_WIDTH  128 
`define AMBA_APB5_USER_DATA_WIDTH `AMBA_APB5_DATA_WIDTH/2

`define AMBA_APB5_COMPLETER0_ADDR_SIZE  32'h0000_1000
`define AMBA_APB5_COMPLETER0_ADDR_START 32'h0000_1000
`define AMBA_APB5_COMPLETER0_ADDR_END   `AMBA_APB5_COMPLETER0_ADDR_START + `AMBA_APB5_COMPLETER0_ADDR_SIZE - 1

`define AMBA_APB5_COMPLETER1_ADDR_SIZE  32'h0000_1000
`define AMBA_APB5_COMPLETER1_ADDR_START 32'h0000_3000
`define AMBA_APB5_COMPLETER1_ADDR_END   `AMBA_APB5_COMPLETER1_ADDR_START + `AMBA_APB5_COMPLETER1_ADDR_SIZE - 1
