`include "uvm_macros.svh"

`include "../test/amba_test_package.sv"

module top;
  import uvm_pkg::*;
  import apb5_environment_package::*;
  import amba_environment_package::*;
  import amba_seq_package::*;
  import amba_test_package::*;
  
  logic clock;
  logic resetn;

  logic [     `AMBA_APB5_ADDR_WIDTH-1:0] paddr;
  logic [                           2:0] pprot;
  logic [                           0:0] pselx;
  logic [                           0:0] penable;
  logic [                           0:0] pwrite;
  logic [     `AMBA_APB5_DATA_WIDTH-1:0] pwdata;
  logic [ (`AMBA_APB5_DATA_WIDTH/8)-1:0] pstrb;

  // source : completer
  logic [                           0:0] pready;
  logic [     `AMBA_APB5_DATA_WIDTH-1:0] prdata;
  logic [                           0:0] pslverr;

  // source : requester
  logic [                           0:0] pwakeup;
  logic [ `AMBA_APB5_USER_REQ_WIDTH-1:0] pauser;

  logic [`AMBA_APB5_USER_DATA_WIDTH-1:0] pwuser;

  // source : completer
  logic [`AMBA_APB5_USER_DATA_WIDTH-1:0] pruser;
  logic [`AMBA_APB5_USER_DATA_WIDTH-1:0] pbuser;

  logic completer0_select, completer1_select;
  
  // Function for address range checking
  function logic addr_in_range(logic [31:0] addr, logic [31:0] range_start, logic [31:0] range_end);
    return (addr >= range_start && addr <= range_end);
  endfunction : addr_in_range

  // Address decoding logic to select the completer
  assign completer0_select = addr_in_range(apb5_requester0_if.paddr, `AMBA_APB5_COMPLETER1_ADDR_START, `AMBA_APB5_COMPLETER1_ADDR_END);
  assign completer1_select = addr_in_range(apb5_requester0_if.paddr, `AMBA_APB5_COMPLETER1_ADDR_START, `AMBA_APB5_COMPLETER1_ADDR_END);

  // apb5_interface #(`AMBA_APB5_ADDR_WIDTH, `AMBA_APB5_DATA_WIDTH, `AMBA_APB5_USER_REQ_WIDTH, `AMBA_APB5_USER_DATA_WIDTH) apb5_requester0_if (clock, resetn);

  // apb5_interface #(`AMBA_APB5_ADDR_WIDTH, `AMBA_APB5_DATA_WIDTH, `AMBA_APB5_USER_REQ_WIDTH, `AMBA_APB5_USER_DATA_WIDTH) apb5_completer0_if (clock, resetn);

  // apb5_interface #(`AMBA_APB5_ADDR_WIDTH, `AMBA_APB5_DATA_WIDTH, `AMBA_APB5_USER_REQ_WIDTH, `AMBA_APB5_USER_DATA_WIDTH) apb5_completer1_if (clock, resetn);

  bind top apb5_interface #(`AMBA_APB5_ADDR_WIDTH, `AMBA_APB5_DATA_WIDTH, `AMBA_APB5_USER_REQ_WIDTH, `AMBA_APB5_USER_DATA_WIDTH) apb5_requester0_if (
    .pclk    ( clock   ),
    .presetn ( resetn  ),
    .paddr   ( paddr   ),
    .pprot   ( pprot   ),
    .pselx   ( pselx   ),
    .penable ( penable ),
    .pwrite  ( pwrite  ),
    .pwdata  ( pwdata  ),
    .pstrb   ( pstrb   ),
    .pready  ( pready  ),
    .prdata  ( prdata  ),
    .pslverr ( pslverr ),
    .pwakeup ( pwakeup ),
    .pauser  ( pauser  ),
    .pwuser  ( pwuser  ),
    .pruser  ( pruser  ),
    .pbuser  ( pbuser  )
  );
  initial begin
    uvm_config_db #(virtual apb5_interface #(`AMBA_APB5_ADDR_WIDTH, `AMBA_APB5_DATA_WIDTH, `AMBA_APB5_USER_REQ_WIDTH, `AMBA_APB5_USER_DATA_WIDTH))::set (null, "*", "apb5_requester0_vif", apb5_requester0_if);
  end

  bind top apb5_interface #(`AMBA_APB5_ADDR_WIDTH, `AMBA_APB5_DATA_WIDTH, `AMBA_APB5_USER_REQ_WIDTH, `AMBA_APB5_USER_DATA_WIDTH) apb5_completer0_if (
    .pclk    ( clock   ),
    .presetn ( resetn  ),
    .paddr   ( paddr   ),
    .pprot   ( pprot   ),
    .pselx   ( pselx   ),
    .penable ( penable ),
    .pwrite  ( pwrite  ),
    .pwdata  ( pwdata  ),
    .pstrb   ( pstrb   ),
    .pready  ( pready  ),
    .prdata  ( prdata  ),
    .pslverr ( pslverr ),
    .pwakeup ( pwakeup ),
    .pauser  ( pauser  ),
    .pwuser  ( pwuser  ),
    .pruser  ( pruser  ),
    .pbuser  ( pbuser  )
  );
  initial begin
    uvm_config_db #(virtual apb5_interface #(`AMBA_APB5_ADDR_WIDTH, `AMBA_APB5_DATA_WIDTH, `AMBA_APB5_USER_REQ_WIDTH, `AMBA_APB5_USER_DATA_WIDTH))::set (null, "*", "apb5_completer0_vif", apb5_completer0_if);
  end

  bind top apb5_interface #(`AMBA_APB5_ADDR_WIDTH, `AMBA_APB5_DATA_WIDTH, `AMBA_APB5_USER_REQ_WIDTH, `AMBA_APB5_USER_DATA_WIDTH) apb5_completer1_if (
    .pclk    ( clock   ),
    .presetn ( resetn  ),
    .paddr   ( paddr   ),
    .pprot   ( pprot   ),
    .pselx   ( pselx   ),
    .penable ( penable ),
    .pwrite  ( pwrite  ),
    .pwdata  ( pwdata  ),
    .pstrb   ( pstrb   ),
    .pready  ( pready  ),
    .prdata  ( prdata  ),
    .pslverr ( pslverr ),
    .pwakeup ( pwakeup ),
    .pauser  ( pauser  ),
    .pwuser  ( pwuser  ),
    .pruser  ( pruser  ),
    .pbuser  ( pbuser  )
  );
  initial begin
    uvm_config_db #(virtual apb5_interface #(`AMBA_APB5_ADDR_WIDTH, `AMBA_APB5_DATA_WIDTH, `AMBA_APB5_USER_REQ_WIDTH, `AMBA_APB5_USER_DATA_WIDTH))::set (null, "*", "apb5_completer1_vif", apb5_completer1_if);
  end


  initial begin
    clock = 0;
    resetn = 0;

    repeat(2) @(posedge clock); 

    resetn = 1;
  end
  
  always #5 clock = !clock;
  
  initial begin
    $dumpfile("dump.vcd"); $dumpvars;
    
    // uvm_config_db #(virtual apb5_interface #(`AMBA_APB5_ADDR_WIDTH, `AMBA_APB5_DATA_WIDTH, `AMBA_APB5_USER_REQ_WIDTH, `AMBA_APB5_USER_DATA_WIDTH))::set (null, "*", "apb5_requester0_vif", apb5_requester0_if);
    // uvm_config_db #(virtual apb5_interface #(`AMBA_APB5_ADDR_WIDTH, `AMBA_APB5_DATA_WIDTH, `AMBA_APB5_USER_REQ_WIDTH, `AMBA_APB5_USER_DATA_WIDTH))::set (null, "*", "apb5_completer0_vif", apb5_completer0_if);
    // uvm_config_db #(virtual apb5_interface #(`AMBA_APB5_ADDR_WIDTH, `AMBA_APB5_DATA_WIDTH, `AMBA_APB5_USER_REQ_WIDTH, `AMBA_APB5_USER_DATA_WIDTH))::set (null, "*", "apb5_completer1_vif", apb5_completer1_if);
    
    uvm_top.finish_on_completion = 1;
    
    run_test("amba_apb5_completer_write_read_test");
  end
endmodule : top
