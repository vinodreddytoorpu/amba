
class apb5_completer_driver #(
  parameter int ADDR_WIDTH      = 32,
  parameter int DATA_WIDTH      = 32,
  parameter int USER_REQ_WIDTH  = 128, 
  parameter int USER_DATA_WIDTH = DATA_WIDTH/2
) extends uvm_driver #(apb5_packet #(ADDR_WIDTH, DATA_WIDTH, USER_REQ_WIDTH, USER_DATA_WIDTH));

  `uvm_component_param_utils(apb5_completer_driver #(ADDR_WIDTH, DATA_WIDTH, USER_REQ_WIDTH, USER_DATA_WIDTH))

  virtual apb5_interface #(ADDR_WIDTH, DATA_WIDTH, USER_REQ_WIDTH, USER_DATA_WIDTH) vif;

  apb5_packet #(ADDR_WIDTH, DATA_WIDTH, USER_REQ_WIDTH, USER_DATA_WIDTH) apb5_pkt;

  apb5_completer_config cfg;

  uvm_component parent_comp;

  extern function new(string name = "apb5_completer_driver", uvm_component parent);
  extern function void build_phase(uvm_phase phase);
  extern function void connect_phase(uvm_phase phase);
  extern task main_phase(uvm_phase phase);
endclass : apb5_completer_driver

function apb5_completer_driver::new(string name = "apb5_completer_driver", uvm_component parent);
  super.new(name, parent);
endfunction : new

function void apb5_completer_driver::build_phase(uvm_phase phase);
  super.build_phase(phase);
  parent_comp = get_parent();
  if(cfg == null) `uvm_fatal(get_name(), $psprintf("apb5_completer_config cfg is null, pass it from parent component %0p", parent_comp.get_name()))
endfunction : build_phase

function void apb5_completer_driver::connect_phase(uvm_phase phase);
  super.connect_phase(phase);
  if(!uvm_config_db #(virtual apb5_interface #(ADDR_WIDTH, DATA_WIDTH, USER_REQ_WIDTH, USER_DATA_WIDTH))::get(this, "*", cfg.vif_path, vif)) `uvm_fatal(get_name(), $psprintf("virtual apb5_interface #(%0d, %0d, %0d, %0d) vif is null, check whether %0s set to config_db::set()", ADDR_WIDTH, DATA_WIDTH, USER_REQ_WIDTH, USER_DATA_WIDTH, cfg.vif_path))
endfunction : connect_phase

task apb5_completer_driver::main_phase(uvm_phase phase);
  super.main_phase(phase);

  fork
    begin
      forever begin
        if(vif.presetn == 1'b0) begin
          vif.pready  <= 1'b1; // default ready
          vif.prdata  <= '0;
          vif.pslverr <= 1'b0;
          vif.pruser  <= '0;
          vif.pbuser  <= '0;
        end
        @(vif.cb_completer); 
      end
    end  
    begin
      forever begin
        apb5_pkt = apb5_packet #(ADDR_WIDTH, DATA_WIDTH, USER_REQ_WIDTH, USER_DATA_WIDTH)::type_id::create("apb5_pkt");
        seq_item_port.get_next_item(apb5_pkt);

        while(1) begin
          if(vif.presetn == 1'b0) @(vif.cb_completer); 
          else break;
        end
        if(vif.pclk == 1'b0) @(posedge vif.pclk); // wait for posedge if clk is low

        vif.pready  <= 1'b1;
        vif.prdata  <= 'hdead_beef;
        vif.pslverr <= 1'b0;
        vif.pruser  <= 1'b0;
        vif.pbuser  <= 1'b0;
        // `uvm_info(get_name(), $sformatf("APB5 Completer Driver APB_ACCESS_PHASE | pready = %0h, pprot = %0h, pselx = %0h, penable = %0h, pwrite = %0h, pwdata = %0h, pstrb = %0h, pwakeup = %0h, pauser = %0h, pwuser = %0h", apb5_pkt.addr, apb5_pkt.prot, 1'b1, 1'b0, apb5_pkt.write, apb5_pkt.wdata, apb5_pkt.strb, apb5_pkt.wakeup, apb5_pkt.auser, apb5_pkt.wuser), UVM_LOW)

        seq_item_port.item_done();
      end
    end  
  join_none
endtask : main_phase
